/*module MEM_WB
(
	input clk,
	//TODO
);

always@(negedge clk)
	begin
	
	end
	
endmodule*/